module fabric (clk, res, in_pins, out_pins, addr, data, wr, cs)

//Clock in configuration data for each pin-mux.
//Config data is simple, the number in the register is
//the physical output pin. 
//always @ ... 

//Generate the required muxes here.
//genvar i ...

endmodule
